//=================================================================================
// MIT License
//
// Copyright (c) 2023 - 2024 Adria Babiano Novella
//
// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:
//
// The above copyright notice and this permission notice shall be included in all
// copies or substantial portions of the Software.
//
// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
// SOFTWARE.
//
// Description    : Arithmetic Logic Unit defines for operations.
// Author         : Adria Babiano
// Created        : Jan 09 2024
//
//=================================================================================

`define ADD 5'h00
`define SUB 5'h01
`define MOD 5'h02
`define NEGA 5'h03
`define INCA 5'h04
`define DECA 5'h05
`define PTA 5'h06
`define ROLA 5'h07
`define RORA 5'h08
`define SHLA 5'h09
`define SHLA2 5'h0a
`define SHLA3 5'h0b
`define SHLA4 5'h0c
`define SHLA5 5'h0d
`define SHLA6 5'h0e
`define SHLA7 5'h0f
`define SHLA8 5'h10
`define SHRA 5'h11
`define SHRA2 5'h12
`define SHRA3 5'h13
`define SHRA4 5'h14
`define SHRA5 5'h15
`define SHRA6 5`h16
`define SHRA7 5'h17
`define SHRA8 5'h18
`define AND 5'h19
`define OR 5'h1a
`define NAND 5'h1b
`define NOR 5'h1c
`define XOR 5'h1d
`define XNOR 5'h1e
`define INVA 5'h1f