//=================================================================================
//
// Description    : Template for description
// Author         : Adria Babiano
// Created        : Dec 30 2023
//
//=================================================================================

package parity_types_pkg;

    typedef enum logic [2:0] {EVEN, ODD, MARK, SPACE, NONE} parity_t;

endpackage
