//=================================================================================
//
// Description    : Template for description
// Author         : Adria Babiano
// Created        : Jan 09 2024
//
//=================================================================================

module 7_seg_hex
	#(
	parameter  = 
	)(
	input logic clk,
	input logic rst_n,
	input logic
	output logic
	);

endmodule
