//=================================================================================
//
// Description    : Template for description
// Author         : Adria Babiano
// Created        : Jan 11 2024
//
//=================================================================================

module one_wire
	#(
	parameter  = 
	)(
	input logic clk,
	input logic rst_n,
	input logic
	output logic
	);

endmodule
