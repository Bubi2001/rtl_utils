`timescale 1ns/1ps

module parity_compute_tb ();
    
endmodule
